../public/chips/C74LS90.vhd