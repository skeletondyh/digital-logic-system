../public/chips/C74LS00.vhd