../public/chips/C74LS20.vhd