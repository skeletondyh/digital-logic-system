../public/chips/C74LS86.vhd