../public/chips/C74LS160.vhd