../public/chips/CD4011.vhd