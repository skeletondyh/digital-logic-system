../public/chips/C74LS27.vhd