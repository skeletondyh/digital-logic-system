../public/chips/C74LS11.vhd