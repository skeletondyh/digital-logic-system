../public/chips/C74LS74.vhd