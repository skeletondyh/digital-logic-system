../public/chips/C74LS14.vhd