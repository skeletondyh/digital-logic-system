../public/chips/C74LS04.vhd