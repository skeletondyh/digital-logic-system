COMPONENT C74LS00 IS 
	PORT (
		port1 : IN  STD_LOGIC;
		port2 : IN  STD_LOGIC;
		port3 : OUT STD_LOGIC;
		port4 : OUT STD_LOGIC;
		port5 : IN  STD_LOGIC;
		port6 : IN  STD_LOGIC;
		port7 : IN  STD_LOGIC; -- GND
		port8 : IN  STD_LOGIC;
		port9 : IN  STD_LOGIC;
		port10: OUT STD_LOGIC;
		port11: OUT STD_LOGIC;
		port12: IN  STD_LOGIC;
		port13: IN  STD_LOGIC;
		port14: IN  STD_LOGIC -- VCC 5V
	);
END C74LS00;