../public/chips/C74LS75.vhd